/* order matters*/
package pck;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "Transaction.svh"
    `include "Sequence.svh"
    `include "Sequencer.svh"
    `include "Driver.svh"
    `include "Monitor.svh"
    `include "Agent.svh"
    `include "Scoreboard.svh"
    `include "Subscriber.svh"
    `include "Env.svh"
    `include "Test.svh"
endpackage